entity mips is
    port 
    (
        clk : in std_logic;
        reset : in std_logic;
    );
end mips;